class home;
  string switch;
  string fan = "OFF";

  extern function void display();
endclass

function void home::display();
  string switch="OFF";
  $display("The switch is %0s that's why fan is %0s",fan,switch);
endfunction:display

module extern_example;
  home h;
  initial begin
    h=new();
    h.display();
  end

endmodule
