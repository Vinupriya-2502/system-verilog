module repeat_code;
initial begin ;
repeat(4)begin  
  $display ("Good morning");
  $display ("Keep shining");
end 
end 
endmodule
