module func_return_void;
  function void display(string str);
    $display("%s",str);
  endfunction 
endmodule 
