interface count_if #(parameter N=4);
  logic rst,clk;
  logic [N:0] counter;
  logic [N:0] counter_up;
endinterface
  
