module top();
  count_if#(2) intf();
  up_counter u1(intf);
  upcounter_testbench u2(intf);
endmodule:top
